entity COMPARATOR_14_BITI_CAT_VREA_CAT_ARE_UTILIZATORUL is
	port
	(
		CAT_VREA,CAT_ARE:in bit_vector(13 downto 0);
		REZULTAT : out bit
	);
end COMPARATOR_14_BITI_CAT_VREA_CAT_ARE_UTILIZATORUL;

architecture AH_COMPARATOR_14_BITI_CAT_VREA_CAT_ARE_UTILIZATORUL of COMPARATOR_14_BITI_CAT_VREA_CAT_ARE_UTILIZATORUL is	
begin
	Comparare:process(CAT_VREA,CAT_ARE)
		begin				 
			if(CAT_VREA<=CAT_ARE) then REZULTAT<='1';
			else REZULTAT<='0';
			end if;
		end process Comparare;
end AH_COMPARATOR_14_BITI_CAT_VREA_CAT_ARE_UTILIZATORUL;